module demultiplexSensor(clk, End, y);
	input clk;
	input [7:0] End;
	output reg [31:0] y;
	
	always @(posedge clk) begin
		case(End)
			8'b00000001: y = 32'b10000000000000000000000000000000;
			8'b00000010: y = 32'b01000000000000000000000000000000;
			8'b00000011: y = 32'b00100000000000000000000000000000;
			8'b00000100: y = 32'b00010000000000000000000000000000;
			8'b00000101: y = 32'b00001000000000000000000000000000;
			8'b00000110: y = 32'b00000100000000000000000000000000;
			8'b00000111: y = 32'b00000010000000000000000000000000;
			8'b00001000: y = 32'b00000001000000000000000000000000;
			8'b00001001: y = 32'b00000000100000000000000000000000;
			8'b00001010: y = 32'b00000000010000000000000000000000;
			8'b00001011: y = 32'b00000000001000000000000000000000;
			8'b00001100: y = 32'b00000000000100000000000000000000;
			8'b00001101: y = 32'b00000000000010000000000000000000;
			8'b00001110: y = 32'b00000000000001000000000000000000;
			8'b00001111: y = 32'b00000000000000100000000000000000;
			8'b00010000: y = 32'b00000000000000010000000000000000;
			8'b00010001: y = 32'b00000000000000001000000000000000;
			8'b00010010: y = 32'b00000000000000000100000000000000;
			8'b00010011: y = 32'b00000000000000000010000000000000;
			8'b00010100: y = 32'b00000000000000000001000000000000;
			8'b00010101: y = 32'b00000000000000000000100000000000;
			8'b00010110: y = 32'b00000000000000000000010000000000;
			8'b00010111: y = 32'b00000000000000000000001000000000;
			8'b00011000: y = 32'b00000000000000000000000100000000;
			8'b00011001: y = 32'b00000000000000000000000010000000;
			8'b00011010: y = 32'b00000000000000000000000001000000;
			8'b00011011: y = 32'b00000000000000000000000000100000;
			8'b00011100: y = 32'b00000000000000000000000000010000;
			8'b00011101: y = 32'b00000000000000000000000000001000;
			8'b00011110: y = 32'b00000000000000000000000000000100;
			8'b00011111: y = 32'b00000000000000000000000000000010;
			8'b00100000: y = 32'b00000000000000000000000000000001;
		endcase
	end
endmodule